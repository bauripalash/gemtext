module main

fn test_version() {
	assert get_version() == '0.0.1'
}
